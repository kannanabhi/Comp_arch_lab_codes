module main_control_pla()
    input [5:0] op;
    output RegDst,ALUsRC,