module bit32_reg(q,d,clk,reset);
    input d,clk,reset;
    output q;

    