module testmux_16;