module testmux_16;
