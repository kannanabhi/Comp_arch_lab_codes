module mux4to1_gate(out,in,sel);
    